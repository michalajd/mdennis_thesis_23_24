
package quickQ_pkg;

    
    // enumerated type for Value Router control signal

    typedef enum logic [2:0] {VR_DEF, VR_ENQ_COMPARE, VR_DEQ_SWAP, VR_LAST, VR_EMPTY, VR_CNT} vrMode_t;    

endpackage