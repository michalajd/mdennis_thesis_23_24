
package quickQ;

    
    // enumerated type for Value Router control signal

    typedef enum {DEF, ENQ_COMPARE, DEQ_SWAP, LAST, EMPTY, CNT} vrMode_t;    

endpackage